-- Ylopoihsh tou Full adder me 2 HA kai mia OR

library ieee;
use ieee.std_logic_1164.all;

entity Full_adder is
Port(
	x, y, z : in std_logic;
	S, Cout : out std_logic
);
end entity Full_adder;

architecture bhv of Full_adder is
begin
	S    <= (x xor y) xor z;
	Cout <= ((x xor y) and z) or (x and y);
end architecture bhv;